`timescale 1ns / 1ps

module mret_adr_sel(
    input logic clk,
    input logic reset_n,
    input logic clear_counter,
    input logic [31:0] current_pc_if1,
    input logic [31:0] current_pc_if2,
    input logic [31:0] current_pc_id,
    input logic [31:0] current_pc_exe,
    input logic [31:0] current_pc_mem_csr,

    output logic [31:0] mepc_adr
    );
    logic [2:0] count_i;
    logic [2:0] count_o;
    logic count_en;
    logic [31:0]mepc_adress_sel[0:5];

    assign count_i = count_o;
    assign count_en = (count_o <=3);

    assign mepc_adress_sel[0] = current_pc_if1;
    assign mepc_adress_sel[1] = current_pc_if2;
    assign mepc_adress_sel[2] = current_pc_id;
    assign mepc_adress_sel[3] = current_pc_exe;
    assign mepc_adress_sel[4] = current_pc_mem_csr;

    n_bit_count_wclr #(.n(3)) counter_reg(
        .clk(clk),
        .reset_n(reset_n),
        .clear(clear_counter),
        .wen(count_en),
        .data_i(count_i),
        .data_o(count_o) );


    assign mepc_adr = mepc_adress_sel[count_o];

//    mux4x1 #(.n(32)) pc_mux(
//        .in0(current_pc_if1),
//        .in1(current_pc_if2),
//        .in2(current_pc_id),
//        .in3(current_pc_exe),
//        .out(mepc_adr),
//        .sel(count_o[1:0])
//        );
endmodule


// counter module
module n_bit_count_wclr #(
    parameter n = 8,
    parameter RESET_VALUE = 0,
    parameter CLR_VALUE = 0
)(
    input logic clk, 
    input logic reset_n,

    input logic wen, 
    input logic  [n-1:0] data_i, 
    output logic [n-1:0] data_o,
    input logic clear
);

    logic [n-1:0] n_bit_reg;
    always_ff @(posedge clk, negedge reset_n) begin 
        if(~reset_n)begin 
            n_bit_reg <= RESET_VALUE;
        end else if (clear) begin
            n_bit_reg <= CLR_VALUE; 
        end else if (wen) begin 
            n_bit_reg <= data_i + 1;
        end
    end

    assign data_o = n_bit_reg;
    
endmodule : n_bit_count_wclr
