module int_pipeline_controller (

    input logic [6:0] opcode_id,
    input logic fun7_5_exe,
    input logic [2:0] fun3_exe,
    fun3_mem,
    input logic zero_mem,
    input logic [1:0] alu_op_exe,
    input logic jump_mem,
    input logic branch_mem,
    input logic mret_type,
    input logic interrupt,
    input logic stall_pipl
    input wire mem_to_reg_exe,
    input wire [4:0] rd_exe,
    // input logic ,


    // output logic []

);



endmodule
